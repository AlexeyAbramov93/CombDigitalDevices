module Main (

input addr

);


endmodule
