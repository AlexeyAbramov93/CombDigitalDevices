// Полный сумматор - логическое устройство с тремя входами и двумя выходами
// для сложения трёх чисел: двух слагаемых a (Ai) и b (Bi) и сигнала переноса из 
// предыдущего разряда c_in (C(i-1)). 
// Результатом сложения являются два числа: сумма по модулю sum и 
// сигнал переноса в следующий разряд c_out (Ci).
// В итоге бит переноса становится старшим битом

module FullAdder (

input a,
input b,

input c_in,

output sum,
output c_out 

);

assign sum = (a^b) ^ c_in;
assign c_out = ((a^b) & c_in) ^ (a&b);

endmodule
