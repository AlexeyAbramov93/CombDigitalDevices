// Шифратор — комбинационное устройство, которое преобразует код из одной (любой) 
// системы счисления в двоичный код. Наибольшее распространение в электронике 
// получили шифраторы, преобразующие позиционный десятичный код, в параллельный двоичный.
// Шифратор используют, например, для перевода десятичных чисел, набранных на
// клавиатуре кнопочного пульта управления, в двоичные числа.

module CD (

//сигнальные входа
input	[7:0] inData,

//выходной двоичный сигнал шифратора
output reg [2:0] outData

);

always @(inData) begin
		case (inData[7:0])	
			8'b00000001 : outData = 3'b000;
			8'b00000010 : outData = 3'b001;
			8'b00000100 : outData = 3'b010;
			8'b00001000 : outData = 3'b011;
			8'b00010000 : outData = 3'b100;
			8'b00100000 : outData = 3'b101;
			8'b01000000 : outData = 3'b110;
			8'b10000000 : outData = 3'b111;			
		endcase	
end
	
endmodule
